module buffer1 (
    input  logic        clk,
    input  logic        rst,
    input  logic        flush,
    input  logic [31:0] pc_in,
    input  logic [31:0] instr_in,
    output logic [31:0] pc_out,
    output logic [31:0] instr_out
);

    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            pc_out    <= 32'b0;
            instr_out <= 32'b0;
        end else if (flush) begin
            pc_out    <= 32'b0;
            instr_out <= 32'b0; // NOP (0x00000000 is often treated as illegal or bubble, essentially NOP here)
        end else begin
            pc_out    <= pc_in;
            instr_out <= instr_in;
        end
    end

endmodule
